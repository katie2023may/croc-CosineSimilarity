/*

This is the Floating Point Arithmetic Unit (acting as an ALU)

*/

`timescale 1 ns / 1 ps

module fpu ();



endmodule