/*

This is the Instruction Memory (control strore) for the microgram

*/


module control_store();



endmodule