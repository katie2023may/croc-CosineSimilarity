/*

This is the Reg File to store intermediate values

*/

module reg_file ();



endmodule