/*

This is the Program Counter (CSAR) module

*/

module pc ();



endmodule