/*

This is the Controller module that generates control signals.

To be connected to datapath.sv inside cosine_sim.sv

*/


module controller ();



endmodule