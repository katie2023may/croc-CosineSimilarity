/*

This is the Datapath module

It connects all of the architetural/state elements of the Cosim microprogram

*/

module datapath();



endmodule