/*

This is the TOP MODULE for the Cosine Similarity Algorithm

Implemented as a Microprogram

Instantiated external Floating Point Arithmetic Unit (FPAU)

*/

`timescale 1 ns / 1 ps

module cosine_sim (
  
);




endmodule